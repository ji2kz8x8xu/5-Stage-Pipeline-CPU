module shifter(dataA, dataB, Signal, dataOut);

  input [31:0] dataA, dataB;
  input [5:0]  Signal;
  
  output [31:0] dataOut;
  
  wire [31:0] w1, w2, w3, w4, w5;
  
  parameter SRL = 6'b000010;

  MUX2_1 s0_mux00 (.sel(dataB[0]), .a(dataA[1]),  .b(dataA[0]), .out(w1[0]));
  MUX2_1 s0_mux01 (.sel(dataB[0]), .a(dataA[2]),  .b(dataA[1]), .out(w1[1]));
  MUX2_1 s0_mux02 (.sel(dataB[0]), .a(dataA[3]),  .b(dataA[2]), .out(w1[2]));
  MUX2_1 s0_mux03 (.sel(dataB[0]), .a(dataA[4]),  .b(dataA[3]), .out(w1[3]));
  MUX2_1 s0_mux04 (.sel(dataB[0]), .a(dataA[5]),  .b(dataA[4]), .out(w1[4]));
  MUX2_1 s0_mux05 (.sel(dataB[0]), .a(dataA[6]),  .b(dataA[5]), .out(w1[5]));
  MUX2_1 s0_mux06 (.sel(dataB[0]), .a(dataA[7]),  .b(dataA[6]), .out(w1[6]));
  MUX2_1 s0_mux07 (.sel(dataB[0]), .a(dataA[8]),  .b(dataA[7]), .out(w1[7]));
  MUX2_1 s0_mux08 (.sel(dataB[0]), .a(dataA[9]),  .b(dataA[8]), .out(w1[8]));
  MUX2_1 s0_mux09 (.sel(dataB[0]), .a(dataA[10]), .b(dataA[9]), .out(w1[9]));
  MUX2_1 s0_mux10 (.sel(dataB[0]), .a(dataA[11]), .b(dataA[10]),.out(w1[10]));
  MUX2_1 s0_mux11 (.sel(dataB[0]), .a(dataA[12]), .b(dataA[11]),.out(w1[11]));
  MUX2_1 s0_mux12 (.sel(dataB[0]), .a(dataA[13]), .b(dataA[12]),.out(w1[12]));
  MUX2_1 s0_mux13 (.sel(dataB[0]), .a(dataA[14]), .b(dataA[13]),.out(w1[13]));
  MUX2_1 s0_mux14 (.sel(dataB[0]), .a(dataA[15]), .b(dataA[14]),.out(w1[14]));
  MUX2_1 s0_mux15 (.sel(dataB[0]), .a(dataA[16]), .b(dataA[15]),.out(w1[15]));
  MUX2_1 s0_mux16 (.sel(dataB[0]), .a(dataA[17]), .b(dataA[16]),.out(w1[16]));
  MUX2_1 s0_mux17 (.sel(dataB[0]), .a(dataA[18]), .b(dataA[17]),.out(w1[17]));
  MUX2_1 s0_mux18 (.sel(dataB[0]), .a(dataA[19]), .b(dataA[18]),.out(w1[18]));
  MUX2_1 s0_mux19 (.sel(dataB[0]), .a(dataA[20]), .b(dataA[19]),.out(w1[19]));
  MUX2_1 s0_mux20 (.sel(dataB[0]), .a(dataA[21]), .b(dataA[20]),.out(w1[20]));
  MUX2_1 s0_mux21 (.sel(dataB[0]), .a(dataA[22]), .b(dataA[21]),.out(w1[21]));
  MUX2_1 s0_mux22 (.sel(dataB[0]), .a(dataA[23]), .b(dataA[22]),.out(w1[22]));
  MUX2_1 s0_mux23 (.sel(dataB[0]), .a(dataA[24]), .b(dataA[23]),.out(w1[23]));
  MUX2_1 s0_mux24 (.sel(dataB[0]), .a(dataA[25]), .b(dataA[24]),.out(w1[24]));
  MUX2_1 s0_mux25 (.sel(dataB[0]), .a(dataA[26]), .b(dataA[25]),.out(w1[25]));
  MUX2_1 s0_mux26 (.sel(dataB[0]), .a(dataA[27]), .b(dataA[26]),.out(w1[26]));
  MUX2_1 s0_mux27 (.sel(dataB[0]), .a(dataA[28]), .b(dataA[27]),.out(w1[27]));
  MUX2_1 s0_mux28 (.sel(dataB[0]), .a(dataA[29]), .b(dataA[28]),.out(w1[28]));
  MUX2_1 s0_mux29 (.sel(dataB[0]), .a(dataA[30]), .b(dataA[29]),.out(w1[29]));
  MUX2_1 s0_mux30 (.sel(dataB[0]), .a(dataA[31]), .b(dataA[30]),.out(w1[30]));
  MUX2_1 s0_mux31 (.sel(dataB[0]), .a(1'b0),      .b(dataA[31]),.out(w1[31]));
  
  MUX2_1 s1_mux00 (.sel(dataB[1]), .a(w1[2]),  .b(w1[0]),  .out(w2[0]));
  MUX2_1 s1_mux01 (.sel(dataB[1]), .a(w1[3]),  .b(w1[1]),  .out(w2[1]));
  MUX2_1 s1_mux02 (.sel(dataB[1]), .a(w1[4]),  .b(w1[2]),  .out(w2[2]));
  MUX2_1 s1_mux03 (.sel(dataB[1]), .a(w1[5]),  .b(w1[3]),  .out(w2[3]));
  MUX2_1 s1_mux04 (.sel(dataB[1]), .a(w1[6]),  .b(w1[4]),  .out(w2[4]));
  MUX2_1 s1_mux05 (.sel(dataB[1]), .a(w1[7]),  .b(w1[5]),  .out(w2[5]));
  MUX2_1 s1_mux06 (.sel(dataB[1]), .a(w1[8]),  .b(w1[6]),  .out(w2[6]));
  MUX2_1 s1_mux07 (.sel(dataB[1]), .a(w1[9]),  .b(w1[7]),  .out(w2[7]));
  MUX2_1 s1_mux08 (.sel(dataB[1]), .a(w1[10]), .b(w1[8]),  .out(w2[8]));
  MUX2_1 s1_mux09 (.sel(dataB[1]), .a(w1[11]), .b(w1[9]),  .out(w2[9]));
  MUX2_1 s1_mux10 (.sel(dataB[1]), .a(w1[12]), .b(w1[10]), .out(w2[10]));
  MUX2_1 s1_mux11 (.sel(dataB[1]), .a(w1[13]), .b(w1[11]), .out(w2[11]));
  MUX2_1 s1_mux12 (.sel(dataB[1]), .a(w1[14]), .b(w1[12]), .out(w2[12]));
  MUX2_1 s1_mux13 (.sel(dataB[1]), .a(w1[15]), .b(w1[13]), .out(w2[13]));
  MUX2_1 s1_mux14 (.sel(dataB[1]), .a(w1[16]), .b(w1[14]), .out(w2[14]));
  MUX2_1 s1_mux15 (.sel(dataB[1]), .a(w1[17]), .b(w1[15]), .out(w2[15]));
  MUX2_1 s1_mux16 (.sel(dataB[1]), .a(w1[18]), .b(w1[16]), .out(w2[16]));
  MUX2_1 s1_mux17 (.sel(dataB[1]), .a(w1[19]), .b(w1[17]), .out(w2[17]));
  MUX2_1 s1_mux18 (.sel(dataB[1]), .a(w1[20]), .b(w1[18]), .out(w2[18]));
  MUX2_1 s1_mux19 (.sel(dataB[1]), .a(w1[21]), .b(w1[19]), .out(w2[19]));
  MUX2_1 s1_mux20 (.sel(dataB[1]), .a(w1[22]), .b(w1[20]), .out(w2[20]));
  MUX2_1 s1_mux21 (.sel(dataB[1]), .a(w1[23]), .b(w1[21]), .out(w2[21]));
  MUX2_1 s1_mux22 (.sel(dataB[1]), .a(w1[24]), .b(w1[22]), .out(w2[22]));
  MUX2_1 s1_mux23 (.sel(dataB[1]), .a(w1[25]), .b(w1[23]), .out(w2[23]));
  MUX2_1 s1_mux24 (.sel(dataB[1]), .a(w1[26]), .b(w1[24]), .out(w2[24]));
  MUX2_1 s1_mux25 (.sel(dataB[1]), .a(w1[27]), .b(w1[25]), .out(w2[25]));
  MUX2_1 s1_mux26 (.sel(dataB[1]), .a(w1[28]), .b(w1[26]), .out(w2[26]));
  MUX2_1 s1_mux27 (.sel(dataB[1]), .a(w1[29]), .b(w1[27]), .out(w2[27]));
  MUX2_1 s1_mux28 (.sel(dataB[1]), .a(w1[30]), .b(w1[28]), .out(w2[28]));
  MUX2_1 s1_mux29 (.sel(dataB[1]), .a(w1[31]), .b(w1[29]), .out(w2[29]));
  MUX2_1 s1_mux30 (.sel(dataB[1]), .a(1'b0),   .b(w1[30]), .out(w2[30]));
  MUX2_1 s1_mux31 (.sel(dataB[1]), .a(1'b0),   .b(w1[31]), .out(w2[31]));

  MUX2_1 s2_mux00 (.sel(dataB[2]), .a(w2[4]),  .b(w2[0]),  .out(w3[0]));
  MUX2_1 s2_mux01 (.sel(dataB[2]), .a(w2[5]),  .b(w2[1]),  .out(w3[1]));
  MUX2_1 s2_mux02 (.sel(dataB[2]), .a(w2[6]),  .b(w2[2]),  .out(w3[2]));
  MUX2_1 s2_mux03 (.sel(dataB[2]), .a(w2[7]),  .b(w2[3]),  .out(w3[3]));
  MUX2_1 s2_mux04 (.sel(dataB[2]), .a(w2[8]),  .b(w2[4]),  .out(w3[4]));
  MUX2_1 s2_mux05 (.sel(dataB[2]), .a(w2[9]),  .b(w2[5]),  .out(w3[5]));
  MUX2_1 s2_mux06 (.sel(dataB[2]), .a(w2[10]), .b(w2[6]),  .out(w3[6]));
  MUX2_1 s2_mux07 (.sel(dataB[2]), .a(w2[11]), .b(w2[7]),  .out(w3[7]));
  MUX2_1 s2_mux08 (.sel(dataB[2]), .a(w2[12]), .b(w2[8]),  .out(w3[8]));
  MUX2_1 s2_mux09 (.sel(dataB[2]), .a(w2[13]), .b(w2[9]),  .out(w3[9]));
  MUX2_1 s2_mux10 (.sel(dataB[2]), .a(w2[14]), .b(w2[10]), .out(w3[10]));
  MUX2_1 s2_mux11 (.sel(dataB[2]), .a(w2[15]), .b(w2[11]), .out(w3[11]));
  MUX2_1 s2_mux12 (.sel(dataB[2]), .a(w2[16]), .b(w2[12]), .out(w3[12]));
  MUX2_1 s2_mux13 (.sel(dataB[2]), .a(w2[17]), .b(w2[13]), .out(w3[13]));
  MUX2_1 s2_mux14 (.sel(dataB[2]), .a(w2[18]), .b(w2[14]), .out(w3[14]));
  MUX2_1 s2_mux15 (.sel(dataB[2]), .a(w2[19]), .b(w2[15]), .out(w3[15]));
  MUX2_1 s2_mux16 (.sel(dataB[2]), .a(w2[20]), .b(w2[16]), .out(w3[16]));
  MUX2_1 s2_mux17 (.sel(dataB[2]), .a(w2[21]), .b(w2[17]), .out(w3[17]));
  MUX2_1 s2_mux18 (.sel(dataB[2]), .a(w2[22]), .b(w2[18]), .out(w3[18]));
  MUX2_1 s2_mux19 (.sel(dataB[2]), .a(w2[23]), .b(w2[19]), .out(w3[19]));
  MUX2_1 s2_mux20 (.sel(dataB[2]), .a(w2[24]), .b(w2[20]), .out(w3[20]));
  MUX2_1 s2_mux21 (.sel(dataB[2]), .a(w2[25]), .b(w2[21]), .out(w3[21]));
  MUX2_1 s2_mux22 (.sel(dataB[2]), .a(w2[26]), .b(w2[22]), .out(w3[22]));
  MUX2_1 s2_mux23 (.sel(dataB[2]), .a(w2[27]), .b(w2[23]), .out(w3[23]));
  MUX2_1 s2_mux24 (.sel(dataB[2]), .a(w2[28]), .b(w2[24]), .out(w3[24]));
  MUX2_1 s2_mux25 (.sel(dataB[2]), .a(w2[29]), .b(w2[25]), .out(w3[25]));
  MUX2_1 s2_mux26 (.sel(dataB[2]), .a(w2[30]), .b(w2[26]), .out(w3[26]));
  MUX2_1 s2_mux27 (.sel(dataB[2]), .a(w2[31]), .b(w2[27]), .out(w3[27]));
  MUX2_1 s2_mux28 (.sel(dataB[2]), .a(1'b0),   .b(w2[28]), .out(w3[28]));
  MUX2_1 s2_mux29 (.sel(dataB[2]), .a(1'b0),   .b(w2[29]), .out(w3[29]));
  MUX2_1 s2_mux30 (.sel(dataB[2]), .a(1'b0),   .b(w2[30]), .out(w3[30]));
  MUX2_1 s2_mux31 (.sel(dataB[2]), .a(1'b0),   .b(w2[31]), .out(w3[31]));

  MUX2_1 s3_mux00 (.sel(dataB[3]), .a(w3[8]),  .b(w3[0]),  .out(w4[0]));
  MUX2_1 s3_mux01 (.sel(dataB[3]), .a(w3[9]),  .b(w3[1]),  .out(w4[1]));
  MUX2_1 s3_mux02 (.sel(dataB[3]), .a(w3[10]), .b(w3[2]),  .out(w4[2]));
  MUX2_1 s3_mux03 (.sel(dataB[3]), .a(w3[11]), .b(w3[3]),  .out(w4[3]));
  MUX2_1 s3_mux04 (.sel(dataB[3]), .a(w3[12]), .b(w3[4]),  .out(w4[4]));
  MUX2_1 s3_mux05 (.sel(dataB[3]), .a(w3[13]), .b(w3[5]),  .out(w4[5]));
  MUX2_1 s3_mux06 (.sel(dataB[3]), .a(w3[14]), .b(w3[6]),  .out(w4[6]));
  MUX2_1 s3_mux07 (.sel(dataB[3]), .a(w3[15]), .b(w3[7]),  .out(w4[7]));
  MUX2_1 s3_mux08 (.sel(dataB[3]), .a(w3[16]), .b(w3[8]),  .out(w4[8]));
  MUX2_1 s3_mux09 (.sel(dataB[3]), .a(w3[17]), .b(w3[9]),  .out(w4[9]));
  MUX2_1 s3_mux10 (.sel(dataB[3]), .a(w3[18]), .b(w3[10]), .out(w4[10]));
  MUX2_1 s3_mux11 (.sel(dataB[3]), .a(w3[19]), .b(w3[11]), .out(w4[11]));
  MUX2_1 s3_mux12 (.sel(dataB[3]), .a(w3[20]), .b(w3[12]), .out(w4[12]));
  MUX2_1 s3_mux13 (.sel(dataB[3]), .a(w3[21]), .b(w3[13]), .out(w4[13]));
  MUX2_1 s3_mux14 (.sel(dataB[3]), .a(w3[22]), .b(w3[14]), .out(w4[14]));
  MUX2_1 s3_mux15 (.sel(dataB[3]), .a(w3[23]), .b(w3[15]), .out(w4[15]));
  MUX2_1 s3_mux16 (.sel(dataB[3]), .a(w3[24]), .b(w3[16]), .out(w4[16]));
  MUX2_1 s3_mux17 (.sel(dataB[3]), .a(w3[25]), .b(w3[17]), .out(w4[17]));
  MUX2_1 s3_mux18 (.sel(dataB[3]), .a(w3[26]), .b(w3[18]), .out(w4[18]));
  MUX2_1 s3_mux19 (.sel(dataB[3]), .a(w3[27]), .b(w3[19]), .out(w4[19]));
  MUX2_1 s3_mux20 (.sel(dataB[3]), .a(w3[28]), .b(w3[20]), .out(w4[20]));
  MUX2_1 s3_mux21 (.sel(dataB[3]), .a(w3[29]), .b(w3[21]), .out(w4[21]));
  MUX2_1 s3_mux22 (.sel(dataB[3]), .a(w3[30]), .b(w3[22]), .out(w4[22]));
  MUX2_1 s3_mux23 (.sel(dataB[3]), .a(w3[31]), .b(w3[23]), .out(w4[23]));
  MUX2_1 s3_mux24 (.sel(dataB[3]), .a(1'b0),   .b(w3[24]), .out(w4[24]));
  MUX2_1 s3_mux25 (.sel(dataB[3]), .a(1'b0),   .b(w3[25]), .out(w4[25]));
  MUX2_1 s3_mux26 (.sel(dataB[3]), .a(1'b0),   .b(w3[26]), .out(w4[26]));
  MUX2_1 s3_mux27 (.sel(dataB[3]), .a(1'b0),   .b(w3[27]), .out(w4[27]));
  MUX2_1 s3_mux28 (.sel(dataB[3]), .a(1'b0),   .b(w3[28]), .out(w4[28]));
  MUX2_1 s3_mux29 (.sel(dataB[3]), .a(1'b0),   .b(w3[29]), .out(w4[29]));
  MUX2_1 s3_mux30 (.sel(dataB[3]), .a(1'b0),   .b(w3[30]), .out(w4[30]));
  MUX2_1 s3_mux31 (.sel(dataB[3]), .a(1'b0),   .b(w3[31]), .out(w4[31]));

  MUX2_1 s4_mux00 (.sel(dataB[4]), .a(w4[16]), .b(w4[0]),  .out(w5[0]));
  MUX2_1 s4_mux01 (.sel(dataB[4]), .a(w4[17]), .b(w4[1]),  .out(w5[1]));
  MUX2_1 s4_mux02 (.sel(dataB[4]), .a(w4[18]), .b(w4[2]),  .out(w5[2]));
  MUX2_1 s4_mux03 (.sel(dataB[4]), .a(w4[19]), .b(w4[3]),  .out(w5[3]));
  MUX2_1 s4_mux04 (.sel(dataB[4]), .a(w4[20]), .b(w4[4]),  .out(w5[4]));
  MUX2_1 s4_mux05 (.sel(dataB[4]), .a(w4[21]), .b(w4[5]),  .out(w5[5]));
  MUX2_1 s4_mux06 (.sel(dataB[4]), .a(w4[22]), .b(w4[6]),  .out(w5[6]));
  MUX2_1 s4_mux07 (.sel(dataB[4]), .a(w4[23]), .b(w4[7]),  .out(w5[7]));
  MUX2_1 s4_mux08 (.sel(dataB[4]), .a(w4[24]), .b(w4[8]),  .out(w5[8]));
  MUX2_1 s4_mux09 (.sel(dataB[4]), .a(w4[25]), .b(w4[9]),  .out(w5[9]));
  MUX2_1 s4_mux10 (.sel(dataB[4]), .a(w4[26]), .b(w4[10]), .out(w5[10]));
  MUX2_1 s4_mux11 (.sel(dataB[4]), .a(w4[27]), .b(w4[11]), .out(w5[11]));
  MUX2_1 s4_mux12 (.sel(dataB[4]), .a(w4[28]), .b(w4[12]), .out(w5[12]));
  MUX2_1 s4_mux13 (.sel(dataB[4]), .a(w4[29]), .b(w4[13]), .out(w5[13]));
  MUX2_1 s4_mux14 (.sel(dataB[4]), .a(w4[30]), .b(w4[14]), .out(w5[14]));
  MUX2_1 s4_mux15 (.sel(dataB[4]), .a(w4[31]), .b(w4[15]), .out(w5[15]));
  MUX2_1 s4_mux16 (.sel(dataB[4]), .a(1'b0),   .b(w4[16]), .out(w5[16]));
  MUX2_1 s4_mux17 (.sel(dataB[4]), .a(1'b0),   .b(w4[17]), .out(w5[17]));
  MUX2_1 s4_mux18 (.sel(dataB[4]), .a(1'b0),   .b(w4[18]), .out(w5[18]));
  MUX2_1 s4_mux19 (.sel(dataB[4]), .a(1'b0),   .b(w4[19]), .out(w5[19]));
  MUX2_1 s4_mux20 (.sel(dataB[4]), .a(1'b0),   .b(w4[20]), .out(w5[20]));
  MUX2_1 s4_mux21 (.sel(dataB[4]), .a(1'b0),   .b(w4[21]), .out(w5[21]));
  MUX2_1 s4_mux22 (.sel(dataB[4]), .a(1'b0),   .b(w4[22]), .out(w5[22]));
  MUX2_1 s4_mux23 (.sel(dataB[4]), .a(1'b0),   .b(w4[23]), .out(w5[23]));
  MUX2_1 s4_mux24 (.sel(dataB[4]), .a(1'b0),   .b(w4[24]), .out(w5[24]));
  MUX2_1 s4_mux25 (.sel(dataB[4]), .a(1'b0),   .b(w4[25]), .out(w5[25]));
  MUX2_1 s4_mux26 (.sel(dataB[4]), .a(1'b0),   .b(w4[26]), .out(w5[26]));
  MUX2_1 s4_mux27 (.sel(dataB[4]), .a(1'b0),   .b(w4[27]), .out(w5[27]));
  MUX2_1 s4_mux28 (.sel(dataB[4]), .a(1'b0),   .b(w4[28]), .out(w5[28]));
  MUX2_1 s4_mux29 (.sel(dataB[4]), .a(1'b0),   .b(w4[29]), .out(w5[29]));
  MUX2_1 s4_mux30 (.sel(dataB[4]), .a(1'b0),   .b(w4[30]), .out(w5[30]));
  MUX2_1 s4_mux31 (.sel(dataB[4]), .a(1'b0),   .b(w4[31]), .out(w5[31]));
  
  // SRL 才輸出 shift 結果
  assign dataOut = (Signal == SRL) ? w5 : dataA;
                  
endmodule